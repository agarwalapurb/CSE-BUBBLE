// Garvit Arora - 200372
// Apurb Agarwal - 200179
module zero(
    input [31:0] a,
    output wire out
);

assign out = (a==0);

endmodule